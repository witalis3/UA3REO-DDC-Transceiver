
module DEBUG2 (
	probe);	

	input	[4:0]	probe;
endmodule
