
module DEBUG (
	probe);	

	input	[47:0]	probe;
endmodule
