
module DEBUG (
	probe);	

	input	[7:0]	probe;
endmodule
