
module DEBUG2 (
	probe);	

	input	[15:0]	probe;
endmodule
