
module DEBUG2 (
	probe);	

	input	[7:0]	probe;
endmodule
