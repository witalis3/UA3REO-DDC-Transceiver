
module DEBUG (
	probe);	

	input	[39:0]	probe;
endmodule
