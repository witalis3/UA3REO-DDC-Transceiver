
module DEBUG (
	probe);	

	input	[61:0]	probe;
endmodule
