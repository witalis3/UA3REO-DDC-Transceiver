// megafunction wizard: %FIR II v18.1%
// GENERATION: XML
// tx_ciccomp.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module tx_ciccomp (
		input  wire        clk,                //                     clk.clk
		input  wire        reset_n,            //                     rst.reset_n
		input  wire [23:0] ast_sink_data,      //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,     //                        .valid
		input  wire [1:0]  ast_sink_error,     //                        .error
		input  wire        ast_sink_sop,       //                        .startofpacket
		input  wire        ast_sink_eop,       //                        .endofpacket
		output wire        ast_sink_ready,     //                        .ready
		output wire [47:0] ast_source_data,    // avalon_streaming_source.data
		output wire        ast_source_valid,   //                        .valid
		output wire [1:0]  ast_source_error,   //                        .error
		input  wire        ast_source_ready,   //                        .ready
		output wire        ast_source_sop,     //                        .startofpacket
		output wire        ast_source_eop,     //                        .endofpacket
		output wire [0:0]  ast_source_channel  //                        .channel
	);

	tx_ciccomp_0002 tx_ciccomp_inst (
		.clk                (clk),                //                     clk.clk
		.reset_n            (reset_n),            //                     rst.reset_n
		.ast_sink_data      (ast_sink_data),      //   avalon_streaming_sink.data
		.ast_sink_valid     (ast_sink_valid),     //                        .valid
		.ast_sink_error     (ast_sink_error),     //                        .error
		.ast_sink_sop       (ast_sink_sop),       //                        .startofpacket
		.ast_sink_eop       (ast_sink_eop),       //                        .endofpacket
		.ast_sink_ready     (ast_sink_ready),     //                        .ready
		.ast_source_data    (ast_source_data),    // avalon_streaming_source.data
		.ast_source_valid   (ast_source_valid),   //                        .valid
		.ast_source_error   (ast_source_error),   //                        .error
		.ast_source_ready   (ast_source_ready),   //                        .ready
		.ast_source_sop     (ast_source_sop),     //                        .startofpacket
		.ast_source_eop     (ast_source_eop),     //                        .endofpacket
		.ast_source_channel (ast_source_channel)  //                        .channel
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2022 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="18.1" >
// Retrieval info: 	<generic name="filterType" value="single" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="symmetryMode" value="sym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="2" />
// Retrieval info: 	<generic name="clockRate" value="187.392" />
// Retrieval info: 	<generic name="clockSlack" value="12" />
// Retrieval info: 	<generic name="inputRate" value="0.048" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="true" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone IV E" />
// Retrieval info: 	<generic name="speedGrade" value="slow" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="100" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="24" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="28.00547,-27.10918,19.6764,-4.287138,-19.57803,51.17325,-88.18962,126.5917,-160.6793,183.3968,-186.9875,163.9278,-108.1903,16.62587,109.5634,-263.6386,432.4929,-596.6616,731.1456,-807.5033,796.8746,-674.2083,422.8634,-39.60776,-461.327,1045.188,-1656.287,2219.912,-2648.109,2848.066,-2734.145,2240.889,-1337.475,39.57715,1580.996,-3393.691,5212.191,-6807.592,7927.899,-8327.308,7797.997,-6206.681,3525.288,141.9622,-4547.702,9302.03,-13896.97,17744.6,-20239.05,20824.77,-19078.76,14781.86,-7986.83,-946.5412,11336.42,-22214.28,32386.77,-40551.03,45424.26,-45910.45,41249.42,-31171.21,15989.91,3331.079,-25211.25,47530.77,-67818.6,83470.09,-92052.65,91587.85,-80868.43,59674.41,-28961.76,-9123.587,51298.45,-93407.2,130739.5,-158539.0,172485.6,-169290.6,147135.8,-106120.4,48415.19,21657.19,-97925.22,172748.3,-237782.6,284718.8,-306310.5,297173.1,-254716.5,179607.7,-76220.2,-47582.82,180725.6,-309943.4,420749.0,-499073.2,532561.7,-512352.7,434111.3,-299329.1,115477.6,103682.6,-339223.8,567902.5,-764537.3,903717.7,-962955.0,924514.3,-778538.5,524056.1,-171261.8,-259125.4,734887.0,-1214971.0,1649588.0,-1984595.0,2161447.0,-2122105.0,1806063.0,-1152833.0,88736.89,1483707.0,-3739434.0,7013818.0,-1.203249E7,1.932583E7,1.932583E7,-1.203249E7,7013818.0,-3739434.0,1483707.0,88736.89,-1152833.0,1806063.0,-2122105.0,2161447.0,-1984595.0,1649588.0,-1214971.0,734887.0,-259125.4,-171261.8,524056.1,-778538.5,924514.3,-962955.0,903717.7,-764537.3,567902.5,-339223.8,103682.6,115477.6,-299329.1,434111.3,-512352.7,532561.7,-499073.2,420749.0,-309943.4,180725.6,-47582.82,-76220.2,179607.7,-254716.5,297173.1,-306310.5,284718.8,-237782.6,172748.3,-97925.22,21657.19,48415.19,-106120.4,147135.8,-169290.6,172485.6,-158539.0,130739.5,-93407.2,51298.45,-9123.587,-28961.76,59674.41,-80868.43,91587.85,-92052.65,83470.09,-67818.6,47530.77,-25211.25,3331.079,15989.91,-31171.21,41249.42,-45910.45,45424.26,-40551.03,32386.77,-22214.28,11336.42,-946.5412,-7986.83,14781.86,-19078.76,20824.77,-20239.05,17744.6,-13896.97,9302.03,-4547.702,141.9622,3525.288,-6206.681,7797.997,-8327.308,7927.899,-6807.592,5212.191,-3393.691,1580.996,39.57715,-1337.475,2240.889,-2734.145,2848.066,-2648.109,2219.912,-1656.287,1045.188,-461.327,-39.60776,422.8634,-674.2083,796.8746,-807.5033,731.1456,-596.6616,432.4929,-263.6386,109.5634,16.62587,-108.1903,163.9278,-186.9875,183.3968,-160.6793,126.5917,-88.18962,51.17325,-19.57803,-4.287138,19.6764,-27.10918,28.00547" />
// Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="16" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffComplex" value="false" />
// Retrieval info: 	<generic name="karatsuba" value="false" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="trunc" />
// Retrieval info: 	<generic name="outMsbBitRem" value="0" />
// Retrieval info: 	<generic name="outLSBRound" value="trunc" />
// Retrieval info: 	<generic name="outLsbBitRem" value="0" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : tx_ciccomp.vo
// RELATED_FILES: tx_ciccomp.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, tx_ciccomp_0002_rtl_core.vhd, tx_ciccomp_0002_ast.vhd, tx_ciccomp_0002.vhd
