
module DEBUG (
	probe);	

	input	[87:0]	probe;
endmodule
