
module DEBUG2 (
	probe);	

	input	[31:0]	probe;
endmodule
